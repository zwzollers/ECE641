module rx #(

) (
    input           i_rx,
    output          o_new,
    output          o_err,
    output [7:0]    o_data
);

endmodule