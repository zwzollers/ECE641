module tx #(

) (
    output          o_rx,
    input           i_start,
    input [7:0]     i_data
);


endmodule